package braminter;
import "BDPI" function Bit#(64) get_rint(Bit#(64) data);


interface Bshifter_IFC;
    method Bit#(64) result(Bit#(64) data);
endinterface

endpackage
